-- Design of registerfile for coefficients

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity registerfilecoe is
  generic(
    constant ROW : natural; -- number of words
   -- constant COL : natural; -- wordlength
    constant NOFW : natural); -- 2^NOFW = Number of words in registerfile
  port (
    readAdd : in std_logic_vector(NOFW-1 downto 0);
    dataOut1 : out std_logic_vector(11 downto 0);
    dataOut2 : out std_logic_vector(11 downto 0));

end entity;

architecture structural of registerfilecoe is

  type registerfile is array (ROW-1 downto 0) of std_logic_vector(11 downto 0); -- registerfile of size ROW x COL
  signal regfileReg1, regfileReg2 : registerfile;

  signal readPtr : unsigned(NOFW-1 downto 0);

begin

    -- address conversion
    readPtr <= (unsigned(readAdd));

    -- output logic
    dataOut1 <= regfileReg1(to_integer(readPtr));
    dataOut2 <= regfileReg2(to_integer(readPtr));

    -- coefficients Real
    regfileReg1(0) <= "011111111111";
    regfileReg1(1) <= "011111111111";
    regfileReg1(2) <= "011111111111";
    regfileReg1(3) <= "011111111111";
    regfileReg1(4) <= "011111111111";
    regfileReg1(5) <= "011111111111";
    regfileReg1(6) <= "011111111111";
    regfileReg1(7) <= "011111111111";
    regfileReg1(8) <= "011111111111";
    regfileReg1(9) <= "011111111111";
    regfileReg1(10) <= "011111111111";
    regfileReg1(11) <= "011111111111";
    regfileReg1(12) <= "011111111111";
    regfileReg1(13) <= "011111111110";
    regfileReg1(14) <= "011111111110";
    regfileReg1(15) <= "011111111110";
    regfileReg1(16) <= "011111111110";
    regfileReg1(17) <= "011111111101";
    regfileReg1(18) <= "011111111101";
    regfileReg1(19) <= "011111111101";
    regfileReg1(20) <= "011111111100";
    regfileReg1(21) <= "011111111100";
    regfileReg1(22) <= "011111111011";
    regfileReg1(23) <= "011111111011";
    regfileReg1(24) <= "011111111010";
    regfileReg1(25) <= "011111111010";
    regfileReg1(26) <= "011111111001";
    regfileReg1(27) <= "011111111001";
    regfileReg1(28) <= "011111111000";
    regfileReg1(29) <= "011111111000";
    regfileReg1(30) <= "011111110111";
    regfileReg1(31) <= "011111110111";
    regfileReg1(32) <= "011111110110";
    regfileReg1(33) <= "011111110110";
    regfileReg1(34) <= "011111110101";
    regfileReg1(35) <= "011111110100";
    regfileReg1(36) <= "011111110100";
    regfileReg1(37) <= "011111110011";
    regfileReg1(38) <= "011111110010";
    regfileReg1(39) <= "011111110001";
    regfileReg1(40) <= "011111110001";
    regfileReg1(41) <= "011111110000";
    regfileReg1(42) <= "011111101111";
    regfileReg1(43) <= "011111101110";
    regfileReg1(44) <= "011111101101";
    regfileReg1(45) <= "011111101101";
    regfileReg1(46) <= "011111101100";
    regfileReg1(47) <= "011111101011";
    regfileReg1(48) <= "011111101010";
    regfileReg1(49) <= "011111101001";
    regfileReg1(50) <= "011111101000";
    regfileReg1(51) <= "011111100111";
    regfileReg1(52) <= "011111100110";
    regfileReg1(53) <= "011111100101";
    regfileReg1(54) <= "011111100100";
    regfileReg1(55) <= "011111100011";
    regfileReg1(56) <= "011111100010";
    regfileReg1(57) <= "011111100001";
    regfileReg1(58) <= "011111100000";
    regfileReg1(59) <= "011111011111";
    regfileReg1(60) <= "011111011101";
    regfileReg1(61) <= "011111011100";
    regfileReg1(62) <= "011111011011";
    regfileReg1(63) <= "011111011010";
    regfileReg1(64) <= "011111011001";
    regfileReg1(65) <= "011111010111";
    regfileReg1(66) <= "011111010110";
    regfileReg1(67) <= "011111010101";
    regfileReg1(68) <= "011111010100";
    regfileReg1(69) <= "011111010010";
    regfileReg1(70) <= "011111010001";
    regfileReg1(71) <= "011111010000";
    regfileReg1(72) <= "011111001110";
    regfileReg1(73) <= "011111001101";
    regfileReg1(74) <= "011111001011";
    regfileReg1(75) <= "011111001010";
    regfileReg1(76) <= "011111001001";
    regfileReg1(77) <= "011111000111";
    regfileReg1(78) <= "011111000110";
    regfileReg1(79) <= "011111000100";
    regfileReg1(80) <= "011111000011";
    regfileReg1(81) <= "011111000001";
    regfileReg1(82) <= "011111000000";
    regfileReg1(83) <= "011110111110";
    regfileReg1(84) <= "011110111100";
    regfileReg1(85) <= "011110111011";
    regfileReg1(86) <= "011110111001";
    regfileReg1(87) <= "011110110111";
    regfileReg1(88) <= "011110110110";
    regfileReg1(89) <= "011110110100";
    regfileReg1(90) <= "011110110010";
    regfileReg1(91) <= "011110110001";
    regfileReg1(92) <= "011110101111";
    regfileReg1(93) <= "011110101101";
    regfileReg1(94) <= "011110101011";
    regfileReg1(95) <= "011110101010";
    regfileReg1(96) <= "011110101000";
    regfileReg1(97) <= "011110100110";
    regfileReg1(98) <= "011110100100";
    regfileReg1(99) <= "011110100010";
    regfileReg1(100) <= "011110100000";
    regfileReg1(101) <= "011110011110";
    regfileReg1(102) <= "011110011101";
    regfileReg1(103) <= "011110011011";
    regfileReg1(104) <= "011110011001";
    regfileReg1(105) <= "011110010111";
    regfileReg1(106) <= "011110010101";
    regfileReg1(107) <= "011110010011";
    regfileReg1(108) <= "011110010001";
    regfileReg1(109) <= "011110001111";
    regfileReg1(110) <= "011110001100";
    regfileReg1(111) <= "011110001010";
    regfileReg1(112) <= "011110001000";
    regfileReg1(113) <= "011110000110";
    regfileReg1(114) <= "011110000100";
    regfileReg1(115) <= "011110000010";
    regfileReg1(116) <= "011110000000";
    regfileReg1(117) <= "011101111101";
    regfileReg1(118) <= "011101111011";
    regfileReg1(119) <= "011101111001";
    regfileReg1(120) <= "011101110111";
    regfileReg1(121) <= "011101110100";
    regfileReg1(122) <= "011101110010";
    regfileReg1(123) <= "011101110000";
    regfileReg1(124) <= "011101101110";
    regfileReg1(125) <= "011101101011";
    regfileReg1(126) <= "011101101001";
    regfileReg1(127) <= "011101100111";
    regfileReg1(128) <= "011101100100";
    regfileReg1(129) <= "011101100010";
    regfileReg1(130) <= "011101011111";
    regfileReg1(131) <= "011101011101";
    regfileReg1(132) <= "011101011010";
    regfileReg1(133) <= "011101011000";
    regfileReg1(134) <= "011101010101";
    regfileReg1(135) <= "011101010011";
    regfileReg1(136) <= "011101010000";
    regfileReg1(137) <= "011101001110";
    regfileReg1(138) <= "011101001011";
    regfileReg1(139) <= "011101001001";
    regfileReg1(140) <= "011101000110";
    regfileReg1(141) <= "011101000011";
    regfileReg1(142) <= "011101000001";
    regfileReg1(143) <= "011100111110";
    regfileReg1(144) <= "011100111011";
    regfileReg1(145) <= "011100111001";
    regfileReg1(146) <= "011100110110";
    regfileReg1(147) <= "011100110011";
    regfileReg1(148) <= "011100110000";
    regfileReg1(149) <= "011100101110";
    regfileReg1(150) <= "011100101011";
    regfileReg1(151) <= "011100101000";
    regfileReg1(152) <= "011100100101";
    regfileReg1(153) <= "011100100010";
    regfileReg1(154) <= "011100100000";
    regfileReg1(155) <= "011100011101";
    regfileReg1(156) <= "011100011010";
    regfileReg1(157) <= "011100010111";
    regfileReg1(158) <= "011100010100";
    regfileReg1(159) <= "011100010001";
    regfileReg1(160) <= "011100001110";
    regfileReg1(161) <= "011100001011";
    regfileReg1(162) <= "011100001000";
    regfileReg1(163) <= "011100000101";
    regfileReg1(164) <= "011100000010";
    regfileReg1(165) <= "011011111111";
    regfileReg1(166) <= "011011111100";
    regfileReg1(167) <= "011011111001";
    regfileReg1(168) <= "011011110110";
    regfileReg1(169) <= "011011110011";
    regfileReg1(170) <= "011011110000";
    regfileReg1(171) <= "011011101101";
    regfileReg1(172) <= "011011101001";
    regfileReg1(173) <= "011011100110";
    regfileReg1(174) <= "011011100011";
    regfileReg1(175) <= "011011100000";
    regfileReg1(176) <= "011011011101";
    regfileReg1(177) <= "011011011001";
    regfileReg1(178) <= "011011010110";
    regfileReg1(179) <= "011011010011";
    regfileReg1(180) <= "011011010000";
    regfileReg1(181) <= "011011001100";
    regfileReg1(182) <= "011011001001";
    regfileReg1(183) <= "011011000110";
    regfileReg1(184) <= "011011000010";
    regfileReg1(185) <= "011010111111";
    regfileReg1(186) <= "011010111100";
    regfileReg1(187) <= "011010111000";
    regfileReg1(188) <= "011010110101";
    regfileReg1(189) <= "011010110001";
    regfileReg1(190) <= "011010101110";
    regfileReg1(191) <= "011010101010";
    regfileReg1(192) <= "011010100111";
    regfileReg1(193) <= "011010100011";
    regfileReg1(194) <= "011010100000";
    regfileReg1(195) <= "011010011100";
    regfileReg1(196) <= "011010011001";
    regfileReg1(197) <= "011010010101";
    regfileReg1(198) <= "011010010010";
    regfileReg1(199) <= "011010001110";
    regfileReg1(200) <= "011010001010";
    regfileReg1(201) <= "011010000111";
    regfileReg1(202) <= "011010000011";
    regfileReg1(203) <= "011001111111";
    regfileReg1(204) <= "011001111100";
    regfileReg1(205) <= "011001111000";
    regfileReg1(206) <= "011001110100";
    regfileReg1(207) <= "011001110001";
    regfileReg1(208) <= "011001101101";
    regfileReg1(209) <= "011001101001";
    regfileReg1(210) <= "011001100101";
    regfileReg1(211) <= "011001100010";
    regfileReg1(212) <= "011001011110";
    regfileReg1(213) <= "011001011010";
    regfileReg1(214) <= "011001010110";
    regfileReg1(215) <= "011001010010";
    regfileReg1(216) <= "011001001111";
    regfileReg1(217) <= "011001001011";
    regfileReg1(218) <= "011001000111";
    regfileReg1(219) <= "011001000011";
    regfileReg1(220) <= "011000111111";
    regfileReg1(221) <= "011000111011";
    regfileReg1(222) <= "011000110111";
    regfileReg1(223) <= "011000110011";
    regfileReg1(224) <= "011000101111";
    regfileReg1(225) <= "011000101011";
    regfileReg1(226) <= "011000100111";
    regfileReg1(227) <= "011000100011";
    regfileReg1(228) <= "011000011111";
    regfileReg1(229) <= "011000011011";
    regfileReg1(230) <= "011000010111";
    regfileReg1(231) <= "011000010011";
    regfileReg1(232) <= "011000001111";
    regfileReg1(233) <= "011000001011";
    regfileReg1(234) <= "011000000111";
    regfileReg1(235) <= "011000000010";
    regfileReg1(236) <= "010111111110";
    regfileReg1(237) <= "010111111010";
    regfileReg1(238) <= "010111110110";
    regfileReg1(239) <= "010111110010";
    regfileReg1(240) <= "010111101101";
    regfileReg1(241) <= "010111101001";
    regfileReg1(242) <= "010111100101";
    regfileReg1(243) <= "010111100001";
    regfileReg1(244) <= "010111011100";
    regfileReg1(245) <= "010111011000";
    regfileReg1(246) <= "010111010100";
    regfileReg1(247) <= "010111010000";
    regfileReg1(248) <= "010111001011";
    regfileReg1(249) <= "010111000111";
    regfileReg1(250) <= "010111000011";
    regfileReg1(251) <= "010110111110";
    regfileReg1(252) <= "010110111010";
    regfileReg1(253) <= "010110110101";
    regfileReg1(254) <= "010110110001";
    regfileReg1(255) <= "010110101101";
    regfileReg1(256) <= "010110101000";



    -- coefficients Imaginary
    regfileReg2(0) <= "000000000000";
    regfileReg2(1) <= "111111111010";
    regfileReg2(2) <= "111111110011";
    regfileReg2(3) <= "111111101101";
    regfileReg2(4) <= "111111100111";
    regfileReg2(5) <= "111111100001";
    regfileReg2(6) <= "111111011010";
    regfileReg2(7) <= "111111010100";
    regfileReg2(8) <= "111111001110";
    regfileReg2(9) <= "111111000111";
    regfileReg2(10) <= "111111000001";
    regfileReg2(11) <= "111110111011";
    regfileReg2(12) <= "111110110101";
    regfileReg2(13) <= "111110101110";
    regfileReg2(14) <= "111110101000";
    regfileReg2(15) <= "111110100010";
    regfileReg2(16) <= "111110011100";
    regfileReg2(17) <= "111110010101";
    regfileReg2(18) <= "111110001111";
    regfileReg2(19) <= "111110001001";
    regfileReg2(20) <= "111110000010";
    regfileReg2(21) <= "111101111100";
    regfileReg2(22) <= "111101110110";
    regfileReg2(23) <= "111101110000";
    regfileReg2(24) <= "111101101001";
    regfileReg2(25) <= "111101100011";
    regfileReg2(26) <= "111101011101";
    regfileReg2(27) <= "111101010111";
    regfileReg2(28) <= "111101010000";
    regfileReg2(29) <= "111101001010";
    regfileReg2(30) <= "111101000100";
    regfileReg2(31) <= "111100111110";
    regfileReg2(32) <= "111100110111";
    regfileReg2(33) <= "111100110001";
    regfileReg2(34) <= "111100101011";
    regfileReg2(35) <= "111100100101";
    regfileReg2(36) <= "111100011110";
    regfileReg2(37) <= "111100011000";
    regfileReg2(38) <= "111100010010";
    regfileReg2(39) <= "111100001100";
    regfileReg2(40) <= "111100000101";
    regfileReg2(41) <= "111011111111";
    regfileReg2(42) <= "111011111001";
    regfileReg2(43) <= "111011110011";
    regfileReg2(44) <= "111011101100";
    regfileReg2(45) <= "111011100110";
    regfileReg2(46) <= "111011100000";
    regfileReg2(47) <= "111011011010";
    regfileReg2(48) <= "111011010011";
    regfileReg2(49) <= "111011001101";
    regfileReg2(50) <= "111011000111";
    regfileReg2(51) <= "111011000001";
    regfileReg2(52) <= "111010111011";
    regfileReg2(53) <= "111010110100";
    regfileReg2(54) <= "111010101110";
    regfileReg2(55) <= "111010101000";
    regfileReg2(56) <= "111010100010";
    regfileReg2(57) <= "111010011100";
    regfileReg2(58) <= "111010010101";
    regfileReg2(59) <= "111010001111";
    regfileReg2(60) <= "111010001001";
    regfileReg2(61) <= "111010000011";
    regfileReg2(62) <= "111001111101";
    regfileReg2(63) <= "111001110111";
    regfileReg2(64) <= "111001110000";
    regfileReg2(65) <= "111001101010";
    regfileReg2(66) <= "111001100100";
    regfileReg2(67) <= "111001011110";
    regfileReg2(68) <= "111001011000";
    regfileReg2(69) <= "111001010010";
    regfileReg2(70) <= "111001001100";
    regfileReg2(71) <= "111001000101";
    regfileReg2(72) <= "111000111111";
    regfileReg2(73) <= "111000111001";
    regfileReg2(74) <= "111000110011";
    regfileReg2(75) <= "111000101101";
    regfileReg2(76) <= "111000100111";
    regfileReg2(77) <= "111000100001";
    regfileReg2(78) <= "111000011011";
    regfileReg2(79) <= "111000010100";
    regfileReg2(80) <= "111000001110";
    regfileReg2(81) <= "111000001000";
    regfileReg2(82) <= "111000000010";
    regfileReg2(83) <= "110111111100";
    regfileReg2(84) <= "110111110110";
    regfileReg2(85) <= "110111110000";
    regfileReg2(86) <= "110111101010";
    regfileReg2(87) <= "110111100100";
    regfileReg2(88) <= "110111011110";
    regfileReg2(89) <= "110111011000";
    regfileReg2(90) <= "110111010010";
    regfileReg2(91) <= "110111001100";
    regfileReg2(92) <= "110111000110";
    regfileReg2(93) <= "110111000000";
    regfileReg2(94) <= "110110111010";
    regfileReg2(95) <= "110110110100";
    regfileReg2(96) <= "110110101101";
    regfileReg2(97) <= "110110100111";
    regfileReg2(98) <= "110110100001";
    regfileReg2(99) <= "110110011011";
    regfileReg2(100) <= "110110010101";
    regfileReg2(101) <= "110110010000";
    regfileReg2(102) <= "110110001010";
    regfileReg2(103) <= "110110000100";
    regfileReg2(104) <= "110101111110";
    regfileReg2(105) <= "110101111000";
    regfileReg2(106) <= "110101110010";
    regfileReg2(107) <= "110101101100";
    regfileReg2(108) <= "110101100110";
    regfileReg2(109) <= "110101100000";
    regfileReg2(110) <= "110101011010";
    regfileReg2(111) <= "110101010100";
    regfileReg2(112) <= "110101001110";
    regfileReg2(113) <= "110101001000";
    regfileReg2(114) <= "110101000010";
    regfileReg2(115) <= "110100111100";
    regfileReg2(116) <= "110100110110";
    regfileReg2(117) <= "110100110001";
    regfileReg2(118) <= "110100101011";
    regfileReg2(119) <= "110100100101";
    regfileReg2(120) <= "110100011111";
    regfileReg2(121) <= "110100011001";
    regfileReg2(122) <= "110100010011";
    regfileReg2(123) <= "110100001101";
    regfileReg2(124) <= "110100001000";
    regfileReg2(125) <= "110100000010";
    regfileReg2(126) <= "110011111100";
    regfileReg2(127) <= "110011110110";
    regfileReg2(128) <= "110011110000";
    regfileReg2(129) <= "110011101010";
    regfileReg2(130) <= "110011100101";
    regfileReg2(131) <= "110011011111";
    regfileReg2(132) <= "110011011001";
    regfileReg2(133) <= "110011010011";
    regfileReg2(134) <= "110011001110";
    regfileReg2(135) <= "110011001000";
    regfileReg2(136) <= "110011000010";
    regfileReg2(137) <= "110010111100";
    regfileReg2(138) <= "110010110111";
    regfileReg2(139) <= "110010110001";
    regfileReg2(140) <= "110010101011";
    regfileReg2(141) <= "110010100101";
    regfileReg2(142) <= "110010100000";
    regfileReg2(143) <= "110010011010";
    regfileReg2(144) <= "110010010100";
    regfileReg2(145) <= "110010001111";
    regfileReg2(146) <= "110010001001";
    regfileReg2(147) <= "110010000011";
    regfileReg2(148) <= "110001111110";
    regfileReg2(149) <= "110001111000";
    regfileReg2(150) <= "110001110010";
    regfileReg2(151) <= "110001101101";
    regfileReg2(152) <= "110001100111";
    regfileReg2(153) <= "110001100010";
    regfileReg2(154) <= "110001011100";
    regfileReg2(155) <= "110001010110";
    regfileReg2(156) <= "110001010001";
    regfileReg2(157) <= "110001001011";
    regfileReg2(158) <= "110001000110";
    regfileReg2(159) <= "110001000000";
    regfileReg2(160) <= "110000111011";
    regfileReg2(161) <= "110000110101";
    regfileReg2(162) <= "110000110000";
    regfileReg2(163) <= "110000101010";
    regfileReg2(164) <= "110000100100";
    regfileReg2(165) <= "110000011111";
    regfileReg2(166) <= "110000011001";
    regfileReg2(167) <= "110000010100";
    regfileReg2(168) <= "110000001111";
    regfileReg2(169) <= "110000001001";
    regfileReg2(170) <= "110000000100";
    regfileReg2(171) <= "101111111110";
    regfileReg2(172) <= "101111111001";
    regfileReg2(173) <= "101111110011";
    regfileReg2(174) <= "101111101110";
    regfileReg2(175) <= "101111101001";
    regfileReg2(176) <= "101111100011";
    regfileReg2(177) <= "101111011110";
    regfileReg2(178) <= "101111011000";
    regfileReg2(179) <= "101111010011";
    regfileReg2(180) <= "101111001110";
    regfileReg2(181) <= "101111001000";
    regfileReg2(182) <= "101111000011";
    regfileReg2(183) <= "101110111110";
    regfileReg2(184) <= "101110111000";
    regfileReg2(185) <= "101110110011";
    regfileReg2(186) <= "101110101110";
    regfileReg2(187) <= "101110101000";
    regfileReg2(188) <= "101110100011";
    regfileReg2(189) <= "101110011110";
    regfileReg2(190) <= "101110011001";
    regfileReg2(191) <= "101110010011";
    regfileReg2(192) <= "101110001110";
    regfileReg2(193) <= "101110001001";
    regfileReg2(194) <= "101110000100";
    regfileReg2(195) <= "101101111111";
    regfileReg2(196) <= "101101111001";
    regfileReg2(197) <= "101101110100";
    regfileReg2(198) <= "101101101111";
    regfileReg2(199) <= "101101101010";
    regfileReg2(200) <= "101101100101";
    regfileReg2(201) <= "101101100000";
    regfileReg2(202) <= "101101011010";
    regfileReg2(203) <= "101101010101";
    regfileReg2(204) <= "101101010000";
    regfileReg2(205) <= "101101001011";
    regfileReg2(206) <= "101101000110";
    regfileReg2(207) <= "101101000001";
    regfileReg2(208) <= "101100111100";
    regfileReg2(209) <= "101100110111";
    regfileReg2(210) <= "101100110010";
    regfileReg2(211) <= "101100101101";
    regfileReg2(212) <= "101100101000";
    regfileReg2(213) <= "101100100011";
    regfileReg2(214) <= "101100011110";
    regfileReg2(215) <= "101100011001";
    regfileReg2(216) <= "101100010100";
    regfileReg2(217) <= "101100001111";
    regfileReg2(218) <= "101100001010";
    regfileReg2(219) <= "101100000101";
    regfileReg2(220) <= "101100000000";
    regfileReg2(221) <= "101011111011";
    regfileReg2(222) <= "101011110111";
    regfileReg2(223) <= "101011110010";
    regfileReg2(224) <= "101011101101";
    regfileReg2(225) <= "101011101000";
    regfileReg2(226) <= "101011100011";
    regfileReg2(227) <= "101011011110";
    regfileReg2(228) <= "101011011001";
    regfileReg2(229) <= "101011010101";
    regfileReg2(230) <= "101011010000";
    regfileReg2(231) <= "101011001011";
    regfileReg2(232) <= "101011000110";
    regfileReg2(233) <= "101011000010";
    regfileReg2(234) <= "101010111101";
    regfileReg2(235) <= "101010111000";
    regfileReg2(236) <= "101010110011";
    regfileReg2(237) <= "101010101111";
    regfileReg2(238) <= "101010101010";
    regfileReg2(239) <= "101010100101";
    regfileReg2(240) <= "101010100001";
    regfileReg2(241) <= "101010011100";
    regfileReg2(242) <= "101010010111";
    regfileReg2(243) <= "101010010011";
    regfileReg2(244) <= "101010001110";
    regfileReg2(245) <= "101010001010";
    regfileReg2(246) <= "101010000101";
    regfileReg2(247) <= "101010000000";
    regfileReg2(248) <= "101001111100";
    regfileReg2(249) <= "101001110111";
    regfileReg2(250) <= "101001110011";
    regfileReg2(251) <= "101001101110";
    regfileReg2(252) <= "101001101010";
    regfileReg2(253) <= "101001100101";
    regfileReg2(254) <= "101001100001";
    regfileReg2(255) <= "101001011100";
    regfileReg2(256) <= "101001011000";


end architecture;
