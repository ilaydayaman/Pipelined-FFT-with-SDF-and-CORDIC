-- Design of registerfile for coefficients

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity coeRegisterfile is
  generic(
    constant ROW : natural; -- number of words
    constant COL : natural; -- wordlength
    constant NOFW : natural); -- 2^NOFW = Number of words in registerfile
  port (
    readAdd1 : in std_logic_vector(NOFW-1 downto 0);
    readAdd2 : in std_logic_vector(NOFW-1 downto 0);
    dataOut1 : out std_logic_vector(COL-1 downto 0);
    dataOut2 : out std_logic_vector(COL-1 downto 0));

end entity;

architecture structural of coeRegisterfile is

  type registerfile is array (ROW-1 downto 0) of std_logic_vector(COL-1 downto 0); -- registerfile of size ROW x COL
  signal regfileReg1, regfileReg2 : registerfile;

  signal readPtr1 : unsigned(NOFW-1 downto 0);
  signal readPtr2 : unsigned(NOFW-1 downto 0);

begin

    -- address conversion
    readPtr1 <= (unsigned(readAdd1));
    readPtr2 <= (unsigned(readAdd2));

    -- output logic
    dataOut1 <= regfileReg1(to_integer(readPtr1));
    dataOut2 <= regfileReg2(to_integer(readPtr2));

    -- coefficients Real
    regfileReg1(0) <= "010000000000";
    regfileReg1(1) <= "010000000000";
    regfileReg1(2) <= "010000000000";
    regfileReg1(3) <= "010000000000";
    regfileReg1(4) <= "010000000000";
    regfileReg1(5) <= "010000000000";
    regfileReg1(6) <= "010000000000";
    regfileReg1(7) <= "010000000000";
    regfileReg1(8) <= "010000000000";
    regfileReg1(9) <= "010000000000";
    regfileReg1(10) <= "010000000000";
    regfileReg1(11) <= "001111111111";
    regfileReg1(12) <= "001111111111";
    regfileReg1(13) <= "001111111111";
    regfileReg1(14) <= "001111111111";
    regfileReg1(15) <= "001111111111";
    regfileReg1(16) <= "001111111111";
    regfileReg1(17) <= "001111111111";
    regfileReg1(18) <= "001111111110";
    regfileReg1(19) <= "001111111110";
    regfileReg1(20) <= "001111111110";
    regfileReg1(21) <= "001111111110";
    regfileReg1(22) <= "001111111110";
    regfileReg1(23) <= "001111111101";
    regfileReg1(24) <= "001111111101";
    regfileReg1(25) <= "001111111101";
    regfileReg1(26) <= "001111111101";
    regfileReg1(27) <= "001111111100";
    regfileReg1(28) <= "001111111100";
    regfileReg1(29) <= "001111111100";
    regfileReg1(30) <= "001111111100";
    regfileReg1(31) <= "001111111011";
    regfileReg1(32) <= "001111111011";
    regfileReg1(33) <= "001111111011";
    regfileReg1(34) <= "001111111010";
    regfileReg1(35) <= "001111111010";
    regfileReg1(36) <= "001111111010";
    regfileReg1(37) <= "001111111001";
    regfileReg1(38) <= "001111111001";
    regfileReg1(39) <= "001111111001";
    regfileReg1(40) <= "001111111000";
    regfileReg1(41) <= "001111111000";
    regfileReg1(42) <= "001111111000";
    regfileReg1(43) <= "001111110111";
    regfileReg1(44) <= "001111110111";
    regfileReg1(45) <= "001111110110";
    regfileReg1(46) <= "001111110110";
    regfileReg1(47) <= "001111110101";
    regfileReg1(48) <= "001111110101";
    regfileReg1(49) <= "001111110100";
    regfileReg1(50) <= "001111110100";
    regfileReg1(51) <= "001111110011";
    regfileReg1(52) <= "001111110011";
    regfileReg1(53) <= "001111110010";
    regfileReg1(54) <= "001111110010";
    regfileReg1(55) <= "001111110001";
    regfileReg1(56) <= "001111110001";
    regfileReg1(57) <= "001111110000";
    regfileReg1(58) <= "001111110000";
    regfileReg1(59) <= "001111101111";
    regfileReg1(60) <= "001111101111";
    regfileReg1(61) <= "001111101110";
    regfileReg1(62) <= "001111101110";
    regfileReg1(63) <= "001111101101";
    regfileReg1(64) <= "001111101100";
    regfileReg1(65) <= "001111101100";
    regfileReg1(66) <= "001111101011";
    regfileReg1(67) <= "001111101010";
    regfileReg1(68) <= "001111101010";
    regfileReg1(69) <= "001111101001";
    regfileReg1(70) <= "001111101000";
    regfileReg1(71) <= "001111101000";
    regfileReg1(72) <= "001111100111";
    regfileReg1(73) <= "001111100110";
    regfileReg1(74) <= "001111100110";
    regfileReg1(75) <= "001111100101";
    regfileReg1(76) <= "001111100100";
    regfileReg1(77) <= "001111100100";
    regfileReg1(78) <= "001111100011";
    regfileReg1(79) <= "001111100010";
    regfileReg1(80) <= "001111100001";
    regfileReg1(81) <= "001111100001";
    regfileReg1(82) <= "001111100000";
    regfileReg1(83) <= "001111011111";
    regfileReg1(84) <= "001111011110";
    regfileReg1(85) <= "001111011101";
    regfileReg1(86) <= "001111011101";
    regfileReg1(87) <= "001111011100";
    regfileReg1(88) <= "001111011011";
    regfileReg1(89) <= "001111011010";
    regfileReg1(90) <= "001111011001";
    regfileReg1(91) <= "001111011000";
    regfileReg1(92) <= "001111010111";
    regfileReg1(93) <= "001111010111";
    regfileReg1(94) <= "001111010110";
    regfileReg1(95) <= "001111010101";
    regfileReg1(96) <= "001111010100";
    regfileReg1(97) <= "001111010011";
    regfileReg1(98) <= "001111010010";
    regfileReg1(99) <= "001111010001";
    regfileReg1(100) <= "001111010000";
    regfileReg1(101) <= "001111001111";
    regfileReg1(102) <= "001111001110";
    regfileReg1(103) <= "001111001101";
    regfileReg1(104) <= "001111001100";
    regfileReg1(105) <= "001111001011";
    regfileReg1(106) <= "001111001010";
    regfileReg1(107) <= "001111001001";
    regfileReg1(108) <= "001111001000";
    regfileReg1(109) <= "001111000111";
    regfileReg1(110) <= "001111000110";
    regfileReg1(111) <= "001111000101";
    regfileReg1(112) <= "001111000100";
    regfileReg1(113) <= "001111000011";
    regfileReg1(114) <= "001111000010";
    regfileReg1(115) <= "001111000001";
    regfileReg1(116) <= "001111000000";
    regfileReg1(117) <= "001110111111";
    regfileReg1(118) <= "001110111110";
    regfileReg1(119) <= "001110111101";
    regfileReg1(120) <= "001110111011";
    regfileReg1(121) <= "001110111010";
    regfileReg1(122) <= "001110111001";
    regfileReg1(123) <= "001110111000";
    regfileReg1(124) <= "001110110111";
    regfileReg1(125) <= "001110110110";
    regfileReg1(126) <= "001110110100";
    regfileReg1(127) <= "001110110011";
    regfileReg1(128) <= "001110110010";
    regfileReg1(129) <= "001110110001";
    regfileReg1(130) <= "001110110000";
    regfileReg1(131) <= "001110101110";
    regfileReg1(132) <= "001110101101";
    regfileReg1(133) <= "001110101100";
    regfileReg1(134) <= "001110101011";
    regfileReg1(135) <= "001110101001";
    regfileReg1(136) <= "001110101000";
    regfileReg1(137) <= "001110100111";
    regfileReg1(138) <= "001110100110";
    regfileReg1(139) <= "001110100100";
    regfileReg1(140) <= "001110100011";
    regfileReg1(141) <= "001110100010";
    regfileReg1(142) <= "001110100000";
    regfileReg1(143) <= "001110011111";
    regfileReg1(144) <= "001110011110";
    regfileReg1(145) <= "001110011100";
    regfileReg1(146) <= "001110011011";
    regfileReg1(147) <= "001110011010";
    regfileReg1(148) <= "001110011000";
    regfileReg1(149) <= "001110010111";
    regfileReg1(150) <= "001110010101";
    regfileReg1(151) <= "001110010100";
    regfileReg1(152) <= "001110010011";
    regfileReg1(153) <= "001110010001";
    regfileReg1(154) <= "001110010000";
    regfileReg1(155) <= "001110001110";
    regfileReg1(156) <= "001110001101";
    regfileReg1(157) <= "001110001011";
    regfileReg1(158) <= "001110001010";
    regfileReg1(159) <= "001110001001";
    regfileReg1(160) <= "001110000111";
    regfileReg1(161) <= "001110000110";
    regfileReg1(162) <= "001110000100";
    regfileReg1(163) <= "001110000011";
    regfileReg1(164) <= "001110000001";
    regfileReg1(165) <= "001110000000";
    regfileReg1(166) <= "001101111110";
    regfileReg1(167) <= "001101111101";
    regfileReg1(168) <= "001101111011";
    regfileReg1(169) <= "001101111001";
    regfileReg1(170) <= "001101111000";
    regfileReg1(171) <= "001101110110";
    regfileReg1(172) <= "001101110101";
    regfileReg1(173) <= "001101110011";
    regfileReg1(174) <= "001101110010";
    regfileReg1(175) <= "001101110000";
    regfileReg1(176) <= "001101101110";
    regfileReg1(177) <= "001101101101";
    regfileReg1(178) <= "001101101011";
    regfileReg1(179) <= "001101101001";
    regfileReg1(180) <= "001101101000";
    regfileReg1(181) <= "001101100110";
    regfileReg1(182) <= "001101100100";
    regfileReg1(183) <= "001101100011";
    regfileReg1(184) <= "001101100001";
    regfileReg1(185) <= "001101011111";
    regfileReg1(186) <= "001101011110";
    regfileReg1(187) <= "001101011100";
    regfileReg1(188) <= "001101011010";
    regfileReg1(189) <= "001101011001";
    regfileReg1(190) <= "001101010111";
    regfileReg1(191) <= "001101010101";
    regfileReg1(192) <= "001101010011";
    regfileReg1(193) <= "001101010010";
    regfileReg1(194) <= "001101010000";
    regfileReg1(195) <= "001101001110";
    regfileReg1(196) <= "001101001100";
    regfileReg1(197) <= "001101001011";
    regfileReg1(198) <= "001101001001";
    regfileReg1(199) <= "001101000111";
    regfileReg1(200) <= "001101000101";
    regfileReg1(201) <= "001101000011";
    regfileReg1(202) <= "001101000010";
    regfileReg1(203) <= "001101000000";
    regfileReg1(204) <= "001100111110";
    regfileReg1(205) <= "001100111100";
    regfileReg1(206) <= "001100111010";
    regfileReg1(207) <= "001100111000";
    regfileReg1(208) <= "001100110110";
    regfileReg1(209) <= "001100110101";
    regfileReg1(210) <= "001100110011";
    regfileReg1(211) <= "001100110001";
    regfileReg1(212) <= "001100101111";
    regfileReg1(213) <= "001100101101";
    regfileReg1(214) <= "001100101011";
    regfileReg1(215) <= "001100101001";
    regfileReg1(216) <= "001100100111";
    regfileReg1(217) <= "001100100101";
    regfileReg1(218) <= "001100100011";
    regfileReg1(219) <= "001100100001";
    regfileReg1(220) <= "001100011111";
    regfileReg1(221) <= "001100011110";
    regfileReg1(222) <= "001100011100";
    regfileReg1(223) <= "001100011010";
    regfileReg1(224) <= "001100011000";
    regfileReg1(225) <= "001100010110";
    regfileReg1(226) <= "001100010100";
    regfileReg1(227) <= "001100010010";
    regfileReg1(228) <= "001100010000";
    regfileReg1(229) <= "001100001110";
    regfileReg1(230) <= "001100001011";
    regfileReg1(231) <= "001100001001";
    regfileReg1(232) <= "001100000111";
    regfileReg1(233) <= "001100000101";
    regfileReg1(234) <= "001100000011";
    regfileReg1(235) <= "001100000001";
    regfileReg1(236) <= "001011111111";
    regfileReg1(237) <= "001011111101";
    regfileReg1(238) <= "001011111011";
    regfileReg1(239) <= "001011111001";
    regfileReg1(240) <= "001011110111";
    regfileReg1(241) <= "001011110101";
    regfileReg1(242) <= "001011110011";
    regfileReg1(243) <= "001011110000";
    regfileReg1(244) <= "001011101110";
    regfileReg1(245) <= "001011101100";
    regfileReg1(246) <= "001011101010";
    regfileReg1(247) <= "001011101000";
    regfileReg1(248) <= "001011100110";
    regfileReg1(249) <= "001011100011";
    regfileReg1(250) <= "001011100001";
    regfileReg1(251) <= "001011011111";
    regfileReg1(252) <= "001011011101";
    regfileReg1(253) <= "001011011011";
    regfileReg1(254) <= "001011011001";
    regfileReg1(255) <= "001011010110";

    -- coefficients Imaginary
    regfileReg2(0) <= "000000000000";
    regfileReg2(1) <= "100000000011";
    regfileReg2(2) <= "100000000110";
    regfileReg2(3) <= "100000001001";
    regfileReg2(4) <= "100000001101";
    regfileReg2(5) <= "100000010000";
    regfileReg2(6) <= "100000010011";
    regfileReg2(7) <= "100000010110";
    regfileReg2(8) <= "100000011001";
    regfileReg2(9) <= "100000011100";
    regfileReg2(10) <= "100000011111";
    regfileReg2(11) <= "100000100011";
    regfileReg2(12) <= "100000100110";
    regfileReg2(13) <= "100000101001";
    regfileReg2(14) <= "100000101100";
    regfileReg2(15) <= "100000101111";
    regfileReg2(16) <= "100000110010";
    regfileReg2(17) <= "100000110101";
    regfileReg2(18) <= "100000111001";
    regfileReg2(19) <= "100000111100";
    regfileReg2(20) <= "100000111111";
    regfileReg2(21) <= "100001000010";
    regfileReg2(22) <= "100001000101";
    regfileReg2(23) <= "100001001000";
    regfileReg2(24) <= "100001001011";
    regfileReg2(25) <= "100001001110";
    regfileReg2(26) <= "100001010010";
    regfileReg2(27) <= "100001010101";
    regfileReg2(28) <= "100001011000";
    regfileReg2(29) <= "100001011011";
    regfileReg2(30) <= "100001011110";
    regfileReg2(31) <= "100001100001";
    regfileReg2(32) <= "100001100100";
    regfileReg2(33) <= "100001100111";
    regfileReg2(34) <= "100001101011";
    regfileReg2(35) <= "100001101110";
    regfileReg2(36) <= "100001110001";
    regfileReg2(37) <= "100001110100";
    regfileReg2(38) <= "100001110111";
    regfileReg2(39) <= "100001111010";
    regfileReg2(40) <= "100001111101";
    regfileReg2(41) <= "100010000000";
    regfileReg2(42) <= "100010000100";
    regfileReg2(43) <= "100010000111";
    regfileReg2(44) <= "100010001010";
    regfileReg2(45) <= "100010001101";
    regfileReg2(46) <= "100010010000";
    regfileReg2(47) <= "100010010011";
    regfileReg2(48) <= "100010010110";
    regfileReg2(49) <= "100010011001";
    regfileReg2(50) <= "100010011100";
    regfileReg2(51) <= "100010100000";
    regfileReg2(52) <= "100010100011";
    regfileReg2(53) <= "100010100110";
    regfileReg2(54) <= "100010101001";
    regfileReg2(55) <= "100010101100";
    regfileReg2(56) <= "100010101111";
    regfileReg2(57) <= "100010110010";
    regfileReg2(58) <= "100010110101";
    regfileReg2(59) <= "100010111000";
    regfileReg2(60) <= "100010111011";
    regfileReg2(61) <= "100010111111";
    regfileReg2(62) <= "100011000010";
    regfileReg2(63) <= "100011000101";
    regfileReg2(64) <= "100011001000";
    regfileReg2(65) <= "100011001011";
    regfileReg2(66) <= "100011001110";
    regfileReg2(67) <= "100011010001";
    regfileReg2(68) <= "100011010100";
    regfileReg2(69) <= "100011010111";
    regfileReg2(70) <= "100011011010";
    regfileReg2(71) <= "100011011101";
    regfileReg2(72) <= "100011100000";
    regfileReg2(73) <= "100011100011";
    regfileReg2(74) <= "100011100110";
    regfileReg2(75) <= "100011101010";
    regfileReg2(76) <= "100011101101";
    regfileReg2(77) <= "100011110000";
    regfileReg2(78) <= "100011110011";
    regfileReg2(79) <= "100011110110";
    regfileReg2(80) <= "100011111001";
    regfileReg2(81) <= "100011111100";
    regfileReg2(82) <= "100011111111";
    regfileReg2(83) <= "100100000010";
    regfileReg2(84) <= "100100000101";
    regfileReg2(85) <= "100100001000";
    regfileReg2(86) <= "100100001011";
    regfileReg2(87) <= "100100001110";
    regfileReg2(88) <= "100100010001";
    regfileReg2(89) <= "100100010100";
    regfileReg2(90) <= "100100010111";
    regfileReg2(91) <= "100100011010";
    regfileReg2(92) <= "100100011101";
    regfileReg2(93) <= "100100100000";
    regfileReg2(94) <= "100100100011";
    regfileReg2(95) <= "100100100110";
    regfileReg2(96) <= "100100101001";
    regfileReg2(97) <= "100100101100";
    regfileReg2(98) <= "100100101111";
    regfileReg2(99) <= "100100110010";
    regfileReg2(100) <= "100100110101";
    regfileReg2(101) <= "100100111000";
    regfileReg2(102) <= "100100111011";
    regfileReg2(103) <= "100100111110";
    regfileReg2(104) <= "100101000001";
    regfileReg2(105) <= "100101000100";
    regfileReg2(106) <= "100101000111";
    regfileReg2(107) <= "100101001010";
    regfileReg2(108) <= "100101001101";
    regfileReg2(109) <= "100101010000";
    regfileReg2(110) <= "100101010011";
    regfileReg2(111) <= "100101010110";
    regfileReg2(112) <= "100101011001";
    regfileReg2(113) <= "100101011100";
    regfileReg2(114) <= "100101011111";
    regfileReg2(115) <= "100101100010";
    regfileReg2(116) <= "100101100101";
    regfileReg2(117) <= "100101101000";
    regfileReg2(118) <= "100101101011";
    regfileReg2(119) <= "100101101110";
    regfileReg2(120) <= "100101110001";
    regfileReg2(121) <= "100101110011";
    regfileReg2(122) <= "100101110110";
    regfileReg2(123) <= "100101111001";
    regfileReg2(124) <= "100101111100";
    regfileReg2(125) <= "100101111111";
    regfileReg2(126) <= "100110000010";
    regfileReg2(127) <= "100110000101";
    regfileReg2(128) <= "100110001000";
    regfileReg2(129) <= "100110001011";
    regfileReg2(130) <= "100110001110";
    regfileReg2(131) <= "100110010001";
    regfileReg2(132) <= "100110010011";
    regfileReg2(133) <= "100110010110";
    regfileReg2(134) <= "100110011001";
    regfileReg2(135) <= "100110011100";
    regfileReg2(136) <= "100110011111";
    regfileReg2(137) <= "100110100010";
    regfileReg2(138) <= "100110100101";
    regfileReg2(139) <= "100110101000";
    regfileReg2(140) <= "100110101010";
    regfileReg2(141) <= "100110101101";
    regfileReg2(142) <= "100110110000";
    regfileReg2(143) <= "100110110011";
    regfileReg2(144) <= "100110110110";
    regfileReg2(145) <= "100110111001";
    regfileReg2(146) <= "100110111011";
    regfileReg2(147) <= "100110111110";
    regfileReg2(148) <= "100111000001";
    regfileReg2(149) <= "100111000100";
    regfileReg2(150) <= "100111000111";
    regfileReg2(151) <= "100111001010";
    regfileReg2(152) <= "100111001100";
    regfileReg2(153) <= "100111001111";
    regfileReg2(154) <= "100111010010";
    regfileReg2(155) <= "100111010101";
    regfileReg2(156) <= "100111011000";
    regfileReg2(157) <= "100111011010";
    regfileReg2(158) <= "100111011101";
    regfileReg2(159) <= "100111100000";
    regfileReg2(160) <= "100111100011";
    regfileReg2(161) <= "100111100101";
    regfileReg2(162) <= "100111101000";
    regfileReg2(163) <= "100111101011";
    regfileReg2(164) <= "100111101110";
    regfileReg2(165) <= "100111110001";
    regfileReg2(166) <= "100111110011";
    regfileReg2(167) <= "100111110110";
    regfileReg2(168) <= "100111111001";
    regfileReg2(169) <= "100111111011";
    regfileReg2(170) <= "100111111110";
    regfileReg2(171) <= "101000000001";
    regfileReg2(172) <= "101000000100";
    regfileReg2(173) <= "101000000110";
    regfileReg2(174) <= "101000001001";
    regfileReg2(175) <= "101000001100";
    regfileReg2(176) <= "101000001110";
    regfileReg2(177) <= "101000010001";
    regfileReg2(178) <= "101000010100";
    regfileReg2(179) <= "101000010111";
    regfileReg2(180) <= "101000011001";
    regfileReg2(181) <= "101000011100";
    regfileReg2(182) <= "101000011111";
    regfileReg2(183) <= "101000100001";
    regfileReg2(184) <= "101000100100";
    regfileReg2(185) <= "101000100110";
    regfileReg2(186) <= "101000101001";
    regfileReg2(187) <= "101000101100";
    regfileReg2(188) <= "101000101110";
    regfileReg2(189) <= "101000110001";
    regfileReg2(190) <= "101000110100";
    regfileReg2(191) <= "101000110110";
    regfileReg2(192) <= "101000111001";
    regfileReg2(193) <= "101000111100";
    regfileReg2(194) <= "101000111110";
    regfileReg2(195) <= "101001000001";
    regfileReg2(196) <= "101001000011";
    regfileReg2(197) <= "101001000110";
    regfileReg2(198) <= "101001001000";
    regfileReg2(199) <= "101001001011";
    regfileReg2(200) <= "101001001110";
    regfileReg2(201) <= "101001010000";
    regfileReg2(202) <= "101001010011";
    regfileReg2(203) <= "101001010101";
    regfileReg2(204) <= "101001011000";
    regfileReg2(205) <= "101001011010";
    regfileReg2(206) <= "101001011101";
    regfileReg2(207) <= "101001011111";
    regfileReg2(208) <= "101001100010";
    regfileReg2(209) <= "101001100101";
    regfileReg2(210) <= "101001100111";
    regfileReg2(211) <= "101001101010";
    regfileReg2(212) <= "101001101100";
    regfileReg2(213) <= "101001101111";
    regfileReg2(214) <= "101001110001";
    regfileReg2(215) <= "101001110100";
    regfileReg2(216) <= "101001110110";
    regfileReg2(217) <= "101001111000";
    regfileReg2(218) <= "101001111011";
    regfileReg2(219) <= "101001111101";
    regfileReg2(220) <= "101010000000";
    regfileReg2(221) <= "101010000010";
    regfileReg2(222) <= "101010000101";
    regfileReg2(223) <= "101010000111";
    regfileReg2(224) <= "101010001010";
    regfileReg2(225) <= "101010001100";
    regfileReg2(226) <= "101010001110";
    regfileReg2(227) <= "101010010001";
    regfileReg2(228) <= "101010010011";
    regfileReg2(229) <= "101010010110";
    regfileReg2(230) <= "101010011000";
    regfileReg2(231) <= "101010011010";
    regfileReg2(232) <= "101010011101";
    regfileReg2(233) <= "101010011111";
    regfileReg2(234) <= "101010100010";
    regfileReg2(235) <= "101010100100";
    regfileReg2(236) <= "101010100110";
    regfileReg2(237) <= "101010101001";
    regfileReg2(238) <= "101010101011";
    regfileReg2(239) <= "101010101101";
    regfileReg2(240) <= "101010110000";
    regfileReg2(241) <= "101010110010";
    regfileReg2(242) <= "101010110100";
    regfileReg2(243) <= "101010110111";
    regfileReg2(244) <= "101010111001";
    regfileReg2(245) <= "101010111011";
    regfileReg2(246) <= "101010111110";
    regfileReg2(247) <= "101011000000";
    regfileReg2(248) <= "101011000010";
    regfileReg2(249) <= "101011000100";
    regfileReg2(250) <= "101011000111";
    regfileReg2(251) <= "101011001001";
    regfileReg2(252) <= "101011001011";
    regfileReg2(253) <= "101011001101";
    regfileReg2(254) <= "101011010000";
    regfileReg2(255) <= "101011010010";

end architecture;
