-- Design of registerfile for coefficients

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity registerfilecoe2 is
  generic(
    constant ROW : natural; -- number of words
   -- constant COL : natural; -- wordlength
    constant NOFW : natural); -- 2^NOFW = Number of words in registerfile
  port (
    readAdd : in std_logic_vector(NOFW-1 downto 0);
    dataOut1 : out std_logic_vector(11 downto 0);
    dataOut2 : out std_logic_vector(11 downto 0));

end registerfilecoe2;

architecture structural of registerfilecoe2 is

  type registerfile is array (ROW-1 downto 0) of std_logic_vector(11 downto 0); -- registerfile of size ROW x COL
  signal regfileReg1, regfileReg2 : registerfile;

  signal readPtr : unsigned(NOFW-1 downto 0);

begin

    -- address conversion
    readPtr <= (unsigned(readAdd));

    -- output logic
    dataOut1 <= regfileReg1(to_integer(readPtr));
    dataOut2 <= regfileReg2(to_integer(readPtr));

    -- coefficients Real
    regfileReg1(0) <= "011111111111";
    regfileReg1(1) <= "011111111111";
    regfileReg1(2) <= "011111111111";
    regfileReg1(3) <= "011111111111";
    regfileReg1(4) <= "011111111111";
    regfileReg1(5) <= "011111111111";
    regfileReg1(6) <= "011111111111";
    regfileReg1(7) <= "011111111110";
    regfileReg1(8) <= "011111111110";
    regfileReg1(9) <= "011111111101";
    regfileReg1(10) <= "011111111100";
    regfileReg1(11) <= "011111111011";
    regfileReg1(12) <= "011111111010";
    regfileReg1(13) <= "011111111001";
    regfileReg1(14) <= "011111111000";
    regfileReg1(15) <= "011111110111";
    regfileReg1(16) <= "011111110110";
    regfileReg1(17) <= "011111110101";
    regfileReg1(18) <= "011111110100";
    regfileReg1(19) <= "011111110010";
    regfileReg1(20) <= "011111110001";
    regfileReg1(21) <= "011111101111";
    regfileReg1(22) <= "011111101101";
    regfileReg1(23) <= "011111101100";
    regfileReg1(24) <= "011111101010";
    regfileReg1(25) <= "011111101000";
    regfileReg1(26) <= "011111100110";
    regfileReg1(27) <= "011111100100";
    regfileReg1(28) <= "011111100010";
    regfileReg1(29) <= "011111100000";
    regfileReg1(30) <= "011111011101";
    regfileReg1(31) <= "011111011011";
    regfileReg1(32) <= "011111011001";
    regfileReg1(33) <= "011111010110";
    regfileReg1(34) <= "011111010100";
    regfileReg1(35) <= "011111010001";
    regfileReg1(36) <= "011111001110";
    regfileReg1(37) <= "011111001011";
    regfileReg1(38) <= "011111001001";
    regfileReg1(39) <= "011111000110";
    regfileReg1(40) <= "011111000011";
    regfileReg1(41) <= "011111000000";
    regfileReg1(42) <= "011110111100";
    regfileReg1(43) <= "011110111001";
    regfileReg1(44) <= "011110110110";
    regfileReg1(45) <= "011110110010";
    regfileReg1(46) <= "011110101111";
    regfileReg1(47) <= "011110101011";
    regfileReg1(48) <= "011110101000";
    regfileReg1(49) <= "011110100100";
    regfileReg1(50) <= "011110100000";
    regfileReg1(51) <= "011110011101";
    regfileReg1(52) <= "011110011001";
    regfileReg1(53) <= "011110010101";
    regfileReg1(54) <= "011110010001";
    regfileReg1(55) <= "011110001100";
    regfileReg1(56) <= "011110001000";
    regfileReg1(57) <= "011110000100";
    regfileReg1(58) <= "011110000000";
    regfileReg1(59) <= "011101111011";
    regfileReg1(60) <= "011101110111";
    regfileReg1(61) <= "011101110010";
    regfileReg1(62) <= "011101101110";
    regfileReg1(63) <= "011101101001";
    regfileReg1(64) <= "011101100100";
    regfileReg1(65) <= "011101011111";
    regfileReg1(66) <= "011101011010";
    regfileReg1(67) <= "011101010101";
    regfileReg1(68) <= "011101010000";
    regfileReg1(69) <= "011101001011";
    regfileReg1(70) <= "011101000110";
    regfileReg1(71) <= "011101000001";
    regfileReg1(72) <= "011100111011";
    regfileReg1(73) <= "011100110110";
    regfileReg1(74) <= "011100110000";
    regfileReg1(75) <= "011100101011";
    regfileReg1(76) <= "011100100101";
    regfileReg1(77) <= "011100100000";
    regfileReg1(78) <= "011100011010";
    regfileReg1(79) <= "011100010100";
    regfileReg1(80) <= "011100001110";
    regfileReg1(81) <= "011100001000";
    regfileReg1(82) <= "011100000010";
    regfileReg1(83) <= "011011111100";
    regfileReg1(84) <= "011011110110";
    regfileReg1(85) <= "011011110000";
    regfileReg1(86) <= "011011101001";
    regfileReg1(87) <= "011011100011";
    regfileReg1(88) <= "011011011101";
    regfileReg1(89) <= "011011010110";
    regfileReg1(90) <= "011011010000";
    regfileReg1(91) <= "011011001001";
    regfileReg1(92) <= "011011000010";
    regfileReg1(93) <= "011010111100";
    regfileReg1(94) <= "011010110101";
    regfileReg1(95) <= "011010101110";
    regfileReg1(96) <= "011010100111";
    regfileReg1(97) <= "011010100000";
    regfileReg1(98) <= "011010011001";
    regfileReg1(99) <= "011010010010";
    regfileReg1(100) <= "011010001010";
    regfileReg1(101) <= "011010000011";
    regfileReg1(102) <= "011001111100";
    regfileReg1(103) <= "011001110100";
    regfileReg1(104) <= "011001101101";
    regfileReg1(105) <= "011001100101";
    regfileReg1(106) <= "011001011110";
    regfileReg1(107) <= "011001010110";
    regfileReg1(108) <= "011001001111";
    regfileReg1(109) <= "011001000111";
    regfileReg1(110) <= "011000111111";
    regfileReg1(111) <= "011000110111";
    regfileReg1(112) <= "011000101111";
    regfileReg1(113) <= "011000100111";
    regfileReg1(114) <= "011000011111";
    regfileReg1(115) <= "011000010111";
    regfileReg1(116) <= "011000001111";
    regfileReg1(117) <= "011000000111";
    regfileReg1(118) <= "010111111110";
    regfileReg1(119) <= "010111110110";
    regfileReg1(120) <= "010111101101";
    regfileReg1(121) <= "010111100101";
    regfileReg1(122) <= "010111011100";
    regfileReg1(123) <= "010111010100";
    regfileReg1(124) <= "010111001011";
    regfileReg1(125) <= "010111000011";
    regfileReg1(126) <= "010110111010";
    regfileReg1(127) <= "010110110001";
    regfileReg1(128) <= "010110101000";


    -- coefficients Imaginary
    regfileReg2(0) <= "000000000000";
    regfileReg2(1) <= "111111110011";
    regfileReg2(2) <= "111111100111";
    regfileReg2(3) <= "111111011010";
    regfileReg2(4) <= "111111001110";
    regfileReg2(5) <= "111111000001";
    regfileReg2(6) <= "111110110101";
    regfileReg2(7) <= "111110101000";
    regfileReg2(8) <= "111110011100";
    regfileReg2(9) <= "111110001111";
    regfileReg2(10) <= "111110000010";
    regfileReg2(11) <= "111101110110";
    regfileReg2(12) <= "111101101001";
    regfileReg2(13) <= "111101011101";
    regfileReg2(14) <= "111101010000";
    regfileReg2(15) <= "111101000100";
    regfileReg2(16) <= "111100110111";
    regfileReg2(17) <= "111100101011";
    regfileReg2(18) <= "111100011110";
    regfileReg2(19) <= "111100010010";
    regfileReg2(20) <= "111100000101";
    regfileReg2(21) <= "111011111001";
    regfileReg2(22) <= "111011101100";
    regfileReg2(23) <= "111011100000";
    regfileReg2(24) <= "111011010011";
    regfileReg2(25) <= "111011000111";
    regfileReg2(26) <= "111010111011";
    regfileReg2(27) <= "111010101110";
    regfileReg2(28) <= "111010100010";
    regfileReg2(29) <= "111010010101";
    regfileReg2(30) <= "111010001001";
    regfileReg2(31) <= "111001111101";
    regfileReg2(32) <= "111001110000";
    regfileReg2(33) <= "111001100100";
    regfileReg2(34) <= "111001011000";
    regfileReg2(35) <= "111001001100";
    regfileReg2(36) <= "111000111111";
    regfileReg2(37) <= "111000110011";
    regfileReg2(38) <= "111000100111";
    regfileReg2(39) <= "111000011011";
    regfileReg2(40) <= "111000001110";
    regfileReg2(41) <= "111000000010";
    regfileReg2(42) <= "110111110110";
    regfileReg2(43) <= "110111101010";
    regfileReg2(44) <= "110111011110";
    regfileReg2(45) <= "110111010010";
    regfileReg2(46) <= "110111000110";
    regfileReg2(47) <= "110110111010";
    regfileReg2(48) <= "110110101101";
    regfileReg2(49) <= "110110100001";
    regfileReg2(50) <= "110110010101";
    regfileReg2(51) <= "110110001010";
    regfileReg2(52) <= "110101111110";
    regfileReg2(53) <= "110101110010";
    regfileReg2(54) <= "110101100110";
    regfileReg2(55) <= "110101011010";
    regfileReg2(56) <= "110101001110";
    regfileReg2(57) <= "110101000010";
    regfileReg2(58) <= "110100110110";
    regfileReg2(59) <= "110100101011";
    regfileReg2(60) <= "110100011111";
    regfileReg2(61) <= "110100010011";
    regfileReg2(62) <= "110100001000";
    regfileReg2(63) <= "110011111100";
    regfileReg2(64) <= "110011110000";
    regfileReg2(65) <= "110011100101";
    regfileReg2(66) <= "110011011001";
    regfileReg2(67) <= "110011001110";
    regfileReg2(68) <= "110011000010";
    regfileReg2(69) <= "110010110111";
    regfileReg2(70) <= "110010101011";
    regfileReg2(71) <= "110010100000";
    regfileReg2(72) <= "110010010100";
    regfileReg2(73) <= "110010001001";
    regfileReg2(74) <= "110001111110";
    regfileReg2(75) <= "110001110010";
    regfileReg2(76) <= "110001100111";
    regfileReg2(77) <= "110001011100";
    regfileReg2(78) <= "110001010001";
    regfileReg2(79) <= "110001000110";
    regfileReg2(80) <= "110000111011";
    regfileReg2(81) <= "110000110000";
    regfileReg2(82) <= "110000100100";
    regfileReg2(83) <= "110000011001";
    regfileReg2(84) <= "110000001111";
    regfileReg2(85) <= "110000000100";
    regfileReg2(86) <= "101111111001";
    regfileReg2(87) <= "101111101110";
    regfileReg2(88) <= "101111100011";
    regfileReg2(89) <= "101111011000";
    regfileReg2(90) <= "101111001110";
    regfileReg2(91) <= "101111000011";
    regfileReg2(92) <= "101110111000";
    regfileReg2(93) <= "101110101110";
    regfileReg2(94) <= "101110100011";
    regfileReg2(95) <= "101110011001";
    regfileReg2(96) <= "101110001110";
    regfileReg2(97) <= "101110000100";
    regfileReg2(98) <= "101101111001";
    regfileReg2(99) <= "101101101111";
    regfileReg2(100) <= "101101100101";
    regfileReg2(101) <= "101101011010";
    regfileReg2(102) <= "101101010000";
    regfileReg2(103) <= "101101000110";
    regfileReg2(104) <= "101100111100";
    regfileReg2(105) <= "101100110010";
    regfileReg2(106) <= "101100101000";
    regfileReg2(107) <= "101100011110";
    regfileReg2(108) <= "101100010100";
    regfileReg2(109) <= "101100001010";
    regfileReg2(110) <= "101100000000";
    regfileReg2(111) <= "101011110111";
    regfileReg2(112) <= "101011101101";
    regfileReg2(113) <= "101011100011";
    regfileReg2(114) <= "101011011001";
    regfileReg2(115) <= "101011010000";
    regfileReg2(116) <= "101011000110";
    regfileReg2(117) <= "101010111101";
    regfileReg2(118) <= "101010110011";
    regfileReg2(119) <= "101010101010";
    regfileReg2(120) <= "101010100001";
    regfileReg2(121) <= "101010010111";
    regfileReg2(122) <= "101010001110";
    regfileReg2(123) <= "101010000101";
    regfileReg2(124) <= "101001111100";
    regfileReg2(125) <= "101001110011";
    regfileReg2(126) <= "101001101010";
    regfileReg2(127) <= "101001100001";
    regfileReg2(128) <= "101001011000";


end architecture;
