-- Design of registerfile for coefficients

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity coeRegisterfile is
  generic(
    constant ROW : natural; -- number of words
    constant COL : natural; -- wordlength
    constant NOFW : natural); -- 2^NOFW = Number of words in registerfile
  port (
    readAdd1 : in std_logic_vector(NOFW-1 downto 0);
    readAdd2 : in std_logic_vector(NOFW-1 downto 0);
    dataOut1 : out std_logic_vector(COL-1 downto 0);
    dataOut2 : out std_logic_vector(COL-1 downto 0));

end entity;

architecture structural of coeRegisterfile is

  type registerfile is array (ROW-1 downto 0) of std_logic_vector(COL-1 downto 0); -- registerfile of size ROW x COL
  signal regfileReg1, regfileReg2 : registerfile;

  signal readPtr1 : unsigned(NOFW-1 downto 0);
  signal readPtr2 : unsigned(NOFW-1 downto 0);

begin

    -- address conversion
    readPtr1 <= (unsigned(readAdd1));
    readPtr2 <= (unsigned(readAdd2));

    -- output logic
    dataOut1 <= regfileReg1(to_integer(readPtr1));
    dataOut2 <= regfileReg2(to_integer(readPtr2));

    -- coefficients Real
    regfileReg1(0) <= "010000000000";
    regfileReg1(1) <= "010000000000";
    regfileReg1(2) <= "010000000000";
    regfileReg1(3) <= "010000000000";
    regfileReg1(4) <= "010000000000";
    regfileReg1(5) <= "010000000000";
    regfileReg1(6) <= "001111111111";
    regfileReg1(7) <= "001111111111";
    regfileReg1(8) <= "001111111111";
    regfileReg1(9) <= "001111111110";
    regfileReg1(10) <= "001111111110";
    regfileReg1(11) <= "001111111110";
    regfileReg1(12) <= "001111111101";
    regfileReg1(13) <= "001111111101";
    regfileReg1(14) <= "001111111100";
    regfileReg1(15) <= "001111111100";
    regfileReg1(16) <= "001111111011";
    regfileReg1(17) <= "001111111010";
    regfileReg1(18) <= "001111111010";
    regfileReg1(19) <= "001111111001";
    regfileReg1(20) <= "001111111000";
    regfileReg1(21) <= "001111111000";
    regfileReg1(22) <= "001111110111";
    regfileReg1(23) <= "001111110110";
    regfileReg1(24) <= "001111110101";
    regfileReg1(25) <= "001111110100";
    regfileReg1(26) <= "001111110011";
    regfileReg1(27) <= "001111110010";
    regfileReg1(28) <= "001111110001";
    regfileReg1(29) <= "001111110000";
    regfileReg1(30) <= "001111101111";
    regfileReg1(31) <= "001111101110";
    regfileReg1(32) <= "001111101100";
    regfileReg1(33) <= "001111101011";
    regfileReg1(34) <= "001111101010";
    regfileReg1(35) <= "001111101000";
    regfileReg1(36) <= "001111100111";
    regfileReg1(37) <= "001111100110";
    regfileReg1(38) <= "001111100100";
    regfileReg1(39) <= "001111100011";
    regfileReg1(40) <= "001111100001";
    regfileReg1(41) <= "001111100000";
    regfileReg1(42) <= "001111011110";
    regfileReg1(43) <= "001111011101";
    regfileReg1(44) <= "001111011011";
    regfileReg1(45) <= "001111011001";
    regfileReg1(46) <= "001111010111";
    regfileReg1(47) <= "001111010110";
    regfileReg1(48) <= "001111010100";
    regfileReg1(49) <= "001111010010";
    regfileReg1(50) <= "001111010000";
    regfileReg1(51) <= "001111001110";
    regfileReg1(52) <= "001111001100";
    regfileReg1(53) <= "001111001010";
    regfileReg1(54) <= "001111001000";
    regfileReg1(55) <= "001111000110";
    regfileReg1(56) <= "001111000100";
    regfileReg1(57) <= "001111000010";
    regfileReg1(58) <= "001111000000";
    regfileReg1(59) <= "001110111110";
    regfileReg1(60) <= "001110111011";
    regfileReg1(61) <= "001110111001";
    regfileReg1(62) <= "001110110111";
    regfileReg1(63) <= "001110110100";
    regfileReg1(64) <= "001110110010";
    regfileReg1(65) <= "001110110000";
    regfileReg1(66) <= "001110101101";
    regfileReg1(67) <= "001110101011";
    regfileReg1(68) <= "001110101000";
    regfileReg1(69) <= "001110100110";
    regfileReg1(70) <= "001110100011";
    regfileReg1(71) <= "001110100000";
    regfileReg1(72) <= "001110011110";
    regfileReg1(73) <= "001110011011";
    regfileReg1(74) <= "001110011000";
    regfileReg1(75) <= "001110010101";
    regfileReg1(76) <= "001110010011";
    regfileReg1(77) <= "001110010000";
    regfileReg1(78) <= "001110001101";
    regfileReg1(79) <= "001110001010";
    regfileReg1(80) <= "001110000111";
    regfileReg1(81) <= "001110000100";
    regfileReg1(82) <= "001110000001";
    regfileReg1(83) <= "001101111110";
    regfileReg1(84) <= "001101111011";
    regfileReg1(85) <= "001101111000";
    regfileReg1(86) <= "001101110101";
    regfileReg1(87) <= "001101110010";
    regfileReg1(88) <= "001101101110";
    regfileReg1(89) <= "001101101011";
    regfileReg1(90) <= "001101101000";
    regfileReg1(91) <= "001101100100";
    regfileReg1(92) <= "001101100001";
    regfileReg1(93) <= "001101011110";
    regfileReg1(94) <= "001101011010";
    regfileReg1(95) <= "001101010111";
    regfileReg1(96) <= "001101010011";
    regfileReg1(97) <= "001101010000";
    regfileReg1(98) <= "001101001100";
    regfileReg1(99) <= "001101001001";
    regfileReg1(100) <= "001101000101";
    regfileReg1(101) <= "001101000010";
    regfileReg1(102) <= "001100111110";
    regfileReg1(103) <= "001100111010";
    regfileReg1(104) <= "001100110110";
    regfileReg1(105) <= "001100110011";
    regfileReg1(106) <= "001100101111";
    regfileReg1(107) <= "001100101011";
    regfileReg1(108) <= "001100100111";
    regfileReg1(109) <= "001100100011";
    regfileReg1(110) <= "001100011111";
    regfileReg1(111) <= "001100011100";
    regfileReg1(112) <= "001100011000";
    regfileReg1(113) <= "001100010100";
    regfileReg1(114) <= "001100010000";
    regfileReg1(115) <= "001100001011";
    regfileReg1(116) <= "001100000111";
    regfileReg1(117) <= "001100000011";
    regfileReg1(118) <= "001011111111";
    regfileReg1(119) <= "001011111011";
    regfileReg1(120) <= "001011110111";
    regfileReg1(121) <= "001011110011";
    regfileReg1(122) <= "001011101110";
    regfileReg1(123) <= "001011101010";
    regfileReg1(124) <= "001011100110";
    regfileReg1(125) <= "001011100001";
    regfileReg1(126) <= "001011011101";
    regfileReg1(127) <= "001011011001";

    -- coefficients Imaginary
    regfileReg2(0) <= "000000000000";
    regfileReg2(1) <= "100000000110";
    regfileReg2(2) <= "100000001101";
    regfileReg2(3) <= "100000010011";
    regfileReg2(4) <= "100000011001";
    regfileReg2(5) <= "100000011111";
    regfileReg2(6) <= "100000100110";
    regfileReg2(7) <= "100000101100";
    regfileReg2(8) <= "100000110010";
    regfileReg2(9) <= "100000111001";
    regfileReg2(10) <= "100000111111";
    regfileReg2(11) <= "100001000101";
    regfileReg2(12) <= "100001001011";
    regfileReg2(13) <= "100001010010";
    regfileReg2(14) <= "100001011000";
    regfileReg2(15) <= "100001011110";
    regfileReg2(16) <= "100001100100";
    regfileReg2(17) <= "100001101011";
    regfileReg2(18) <= "100001110001";
    regfileReg2(19) <= "100001110111";
    regfileReg2(20) <= "100001111101";
    regfileReg2(21) <= "100010000100";
    regfileReg2(22) <= "100010001010";
    regfileReg2(23) <= "100010010000";
    regfileReg2(24) <= "100010010110";
    regfileReg2(25) <= "100010011100";
    regfileReg2(26) <= "100010100011";
    regfileReg2(27) <= "100010101001";
    regfileReg2(28) <= "100010101111";
    regfileReg2(29) <= "100010110101";
    regfileReg2(30) <= "100010111011";
    regfileReg2(31) <= "100011000010";
    regfileReg2(32) <= "100011001000";
    regfileReg2(33) <= "100011001110";
    regfileReg2(34) <= "100011010100";
    regfileReg2(35) <= "100011011010";
    regfileReg2(36) <= "100011100000";
    regfileReg2(37) <= "100011100110";
    regfileReg2(38) <= "100011101101";
    regfileReg2(39) <= "100011110011";
    regfileReg2(40) <= "100011111001";
    regfileReg2(41) <= "100011111111";
    regfileReg2(42) <= "100100000101";
    regfileReg2(43) <= "100100001011";
    regfileReg2(44) <= "100100010001";
    regfileReg2(45) <= "100100010111";
    regfileReg2(46) <= "100100011101";
    regfileReg2(47) <= "100100100011";
    regfileReg2(48) <= "100100101001";
    regfileReg2(49) <= "100100101111";
    regfileReg2(50) <= "100100110101";
    regfileReg2(51) <= "100100111011";
    regfileReg2(52) <= "100101000001";
    regfileReg2(53) <= "100101000111";
    regfileReg2(54) <= "100101001101";
    regfileReg2(55) <= "100101010011";
    regfileReg2(56) <= "100101011001";
    regfileReg2(57) <= "100101011111";
    regfileReg2(58) <= "100101100101";
    regfileReg2(59) <= "100101101011";
    regfileReg2(60) <= "100101110001";
    regfileReg2(61) <= "100101110110";
    regfileReg2(62) <= "100101111100";
    regfileReg2(63) <= "100110000010";
    regfileReg2(64) <= "100110001000";
    regfileReg2(65) <= "100110001110";
    regfileReg2(66) <= "100110010011";
    regfileReg2(67) <= "100110011001";
    regfileReg2(68) <= "100110011111";
    regfileReg2(69) <= "100110100101";
    regfileReg2(70) <= "100110101010";
    regfileReg2(71) <= "100110110000";
    regfileReg2(72) <= "100110110110";
    regfileReg2(73) <= "100110111011";
    regfileReg2(74) <= "100111000001";
    regfileReg2(75) <= "100111000111";
    regfileReg2(76) <= "100111001100";
    regfileReg2(77) <= "100111010010";
    regfileReg2(78) <= "100111011000";
    regfileReg2(79) <= "100111011101";
    regfileReg2(80) <= "100111100011";
    regfileReg2(81) <= "100111101000";
    regfileReg2(82) <= "100111101110";
    regfileReg2(83) <= "100111110011";
    regfileReg2(84) <= "100111111001";
    regfileReg2(85) <= "100111111110";
    regfileReg2(86) <= "101000000100";
    regfileReg2(87) <= "101000001001";
    regfileReg2(88) <= "101000001110";
    regfileReg2(89) <= "101000010100";
    regfileReg2(90) <= "101000011001";
    regfileReg2(91) <= "101000011111";
    regfileReg2(92) <= "101000100100";
    regfileReg2(93) <= "101000101001";
    regfileReg2(94) <= "101000101110";
    regfileReg2(95) <= "101000110100";
    regfileReg2(96) <= "101000111001";
    regfileReg2(97) <= "101000111110";
    regfileReg2(98) <= "101001000011";
    regfileReg2(99) <= "101001001000";
    regfileReg2(100) <= "101001001110";
    regfileReg2(101) <= "101001010011";
    regfileReg2(102) <= "101001011000";
    regfileReg2(103) <= "101001011101";
    regfileReg2(104) <= "101001100010";
    regfileReg2(105) <= "101001100111";
    regfileReg2(106) <= "101001101100";
    regfileReg2(107) <= "101001110001";
    regfileReg2(108) <= "101001110110";
    regfileReg2(109) <= "101001111011";
    regfileReg2(110) <= "101010000000";
    regfileReg2(111) <= "101010000101";
    regfileReg2(112) <= "101010001010";
    regfileReg2(113) <= "101010001110";
    regfileReg2(114) <= "101010010011";
    regfileReg2(115) <= "101010011000";
    regfileReg2(116) <= "101010011101";
    regfileReg2(117) <= "101010100010";
    regfileReg2(118) <= "101010100110";
    regfileReg2(119) <= "101010101011";
    regfileReg2(120) <= "101010110000";
    regfileReg2(121) <= "101010110100";
    regfileReg2(122) <= "101010111001";
    regfileReg2(123) <= "101010111110";
    regfileReg2(124) <= "101011000010";
    regfileReg2(125) <= "101011000111";
    regfileReg2(126) <= "101011001011";
    regfileReg2(127) <= "101011010000";

end architecture;
