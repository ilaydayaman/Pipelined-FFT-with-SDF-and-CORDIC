-- Design of registerfile for coefficients
library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity registerfilecoe2 is
  generic(
    constant ROW  : natural;            -- number of words
    constant NOFW : natural);  -- 2^NOFW = Number of words in registerfile
  port (
    readAdd  : in  std_logic_vector(NOFW-1 downto 0);
    dataOut1 : out std_logic_vector(11 downto 0);
    dataOut2 : out std_logic_vector(11 downto 0));

end registerfilecoe2;

architecture structural of registerfilecoe2 is

  -- registerfile of size ROW x COL
  type registerfile is array (ROW-1 downto 0) of std_logic_vector(11 downto 0);
  signal regfileReg1, regfileReg2 : registerfile;

  signal readPtr : unsigned(NOFW-1 downto 0);

begin

  -- address conversion
  readPtr <= (unsigned(readAdd));

  -- output logic
  dataOut1 <= regfileReg1(to_integer(readPtr));
  dataOut2 <= regfileReg2(to_integer(readPtr));

  -- coefficients Real
  regfileReg1(0)   <= "010000000000";
  regfileReg1(1)   <= "010000000000";
  regfileReg1(2)   <= "010000000000";
  regfileReg1(3)   <= "010000000000";
  regfileReg1(4)   <= "010000000000";
  regfileReg1(5)   <= "010000000000";
  regfileReg1(6)   <= "001111111111";
  regfileReg1(7)   <= "001111111111";
  regfileReg1(8)   <= "001111111111";
  regfileReg1(9)   <= "001111111110";
  regfileReg1(10)  <= "001111111110";
  regfileReg1(11)  <= "001111111110";
  regfileReg1(12)  <= "001111111101";
  regfileReg1(13)  <= "001111111101";
  regfileReg1(14)  <= "001111111100";
  regfileReg1(15)  <= "001111111100";
  regfileReg1(16)  <= "001111111011";
  regfileReg1(17)  <= "001111111010";
  regfileReg1(18)  <= "001111111010";
  regfileReg1(19)  <= "001111111001";
  regfileReg1(20)  <= "001111111000";
  regfileReg1(21)  <= "001111111000";
  regfileReg1(22)  <= "001111110111";
  regfileReg1(23)  <= "001111110110";
  regfileReg1(24)  <= "001111110101";
  regfileReg1(25)  <= "001111110100";
  regfileReg1(26)  <= "001111110011";
  regfileReg1(27)  <= "001111110010";
  regfileReg1(28)  <= "001111110001";
  regfileReg1(29)  <= "001111110000";
  regfileReg1(30)  <= "001111101111";
  regfileReg1(31)  <= "001111101110";
  regfileReg1(32)  <= "001111101100";
  regfileReg1(33)  <= "001111101011";
  regfileReg1(34)  <= "001111101010";
  regfileReg1(35)  <= "001111101000";
  regfileReg1(36)  <= "001111100111";
  regfileReg1(37)  <= "001111100110";
  regfileReg1(38)  <= "001111100100";
  regfileReg1(39)  <= "001111100011";
  regfileReg1(40)  <= "001111100001";
  regfileReg1(41)  <= "001111100000";
  regfileReg1(42)  <= "001111011110";
  regfileReg1(43)  <= "001111011101";
  regfileReg1(44)  <= "001111011011";
  regfileReg1(45)  <= "001111011001";
  regfileReg1(46)  <= "001111010111";
  regfileReg1(47)  <= "001111010110";
  regfileReg1(48)  <= "001111010100";
  regfileReg1(49)  <= "001111010010";
  regfileReg1(50)  <= "001111010000";
  regfileReg1(51)  <= "001111001110";
  regfileReg1(52)  <= "001111001100";
  regfileReg1(53)  <= "001111001010";
  regfileReg1(54)  <= "001111001000";
  regfileReg1(55)  <= "001111000110";
  regfileReg1(56)  <= "001111000100";
  regfileReg1(57)  <= "001111000010";
  regfileReg1(58)  <= "001111000000";
  regfileReg1(59)  <= "001110111110";
  regfileReg1(60)  <= "001110111011";
  regfileReg1(61)  <= "001110111001";
  regfileReg1(62)  <= "001110110111";
  regfileReg1(63)  <= "001110110100";
  regfileReg1(64)  <= "001110110010";
  regfileReg1(65)  <= "001110110000";
  regfileReg1(66)  <= "001110101101";
  regfileReg1(67)  <= "001110101011";
  regfileReg1(68)  <= "001110101000";
  regfileReg1(69)  <= "001110100110";
  regfileReg1(70)  <= "001110100011";
  regfileReg1(71)  <= "001110100000";
  regfileReg1(72)  <= "001110011110";
  regfileReg1(73)  <= "001110011011";
  regfileReg1(74)  <= "001110011000";
  regfileReg1(75)  <= "001110010101";
  regfileReg1(76)  <= "001110010011";
  regfileReg1(77)  <= "001110010000";
  regfileReg1(78)  <= "001110001101";
  regfileReg1(79)  <= "001110001010";
  regfileReg1(80)  <= "001110000111";
  regfileReg1(81)  <= "001110000100";
  regfileReg1(82)  <= "001110000001";
  regfileReg1(83)  <= "001101111110";
  regfileReg1(84)  <= "001101111011";
  regfileReg1(85)  <= "001101111000";
  regfileReg1(86)  <= "001101110101";
  regfileReg1(87)  <= "001101110010";
  regfileReg1(88)  <= "001101101110";
  regfileReg1(89)  <= "001101101011";
  regfileReg1(90)  <= "001101101000";
  regfileReg1(91)  <= "001101100100";
  regfileReg1(92)  <= "001101100001";
  regfileReg1(93)  <= "001101011110";
  regfileReg1(94)  <= "001101011010";
  regfileReg1(95)  <= "001101010111";
  regfileReg1(96)  <= "001101010011";
  regfileReg1(97)  <= "001101010000";
  regfileReg1(98)  <= "001101001100";
  regfileReg1(99)  <= "001101001001";
  regfileReg1(100) <= "001101000101";
  regfileReg1(101) <= "001101000010";
  regfileReg1(102) <= "001100111110";
  regfileReg1(103) <= "001100111010";
  regfileReg1(104) <= "001100110110";
  regfileReg1(105) <= "001100110011";
  regfileReg1(106) <= "001100101111";
  regfileReg1(107) <= "001100101011";
  regfileReg1(108) <= "001100100111";
  regfileReg1(109) <= "001100100011";
  regfileReg1(110) <= "001100011111";
  regfileReg1(111) <= "001100011100";
  regfileReg1(112) <= "001100011000";
  regfileReg1(113) <= "001100010100";
  regfileReg1(114) <= "001100010000";
  regfileReg1(115) <= "001100001011";
  regfileReg1(116) <= "001100000111";
  regfileReg1(117) <= "001100000011";
  regfileReg1(118) <= "001011111111";
  regfileReg1(119) <= "001011111011";
  regfileReg1(120) <= "001011110111";
  regfileReg1(121) <= "001011110011";
  regfileReg1(122) <= "001011101110";
  regfileReg1(123) <= "001011101010";
  regfileReg1(124) <= "001011100110";
  regfileReg1(125) <= "001011100001";
  regfileReg1(126) <= "001011011101";
  regfileReg1(127) <= "001011011001";
  regfileReg1(128) <= "001011010100";

  -- coefficients Imaginary
  regfileReg2(0)   <= "000000000000";
  regfileReg2(1)   <= "111111111010";
  regfileReg2(2)   <= "111111110011";
  regfileReg2(3)   <= "111111101101";
  regfileReg2(4)   <= "111111100111";
  regfileReg2(5)   <= "111111100001";
  regfileReg2(6)   <= "111111011010";
  regfileReg2(7)   <= "111111010100";
  regfileReg2(8)   <= "111111001110";
  regfileReg2(9)   <= "111111000111";
  regfileReg2(10)  <= "111111000001";
  regfileReg2(11)  <= "111110111011";
  regfileReg2(12)  <= "111110110101";
  regfileReg2(13)  <= "111110101110";
  regfileReg2(14)  <= "111110101000";
  regfileReg2(15)  <= "111110100010";
  regfileReg2(16)  <= "111110011100";
  regfileReg2(17)  <= "111110010101";
  regfileReg2(18)  <= "111110001111";
  regfileReg2(19)  <= "111110001001";
  regfileReg2(20)  <= "111110000011";
  regfileReg2(21)  <= "111101111100";
  regfileReg2(22)  <= "111101110110";
  regfileReg2(23)  <= "111101110000";
  regfileReg2(24)  <= "111101101010";
  regfileReg2(25)  <= "111101100100";
  regfileReg2(26)  <= "111101011101";
  regfileReg2(27)  <= "111101010111";
  regfileReg2(28)  <= "111101010001";
  regfileReg2(29)  <= "111101001011";
  regfileReg2(30)  <= "111101000101";
  regfileReg2(31)  <= "111100111110";
  regfileReg2(32)  <= "111100111000";
  regfileReg2(33)  <= "111100110010";
  regfileReg2(34)  <= "111100101100";
  regfileReg2(35)  <= "111100100110";
  regfileReg2(36)  <= "111100100000";
  regfileReg2(37)  <= "111100011010";
  regfileReg2(38)  <= "111100010011";
  regfileReg2(39)  <= "111100001101";
  regfileReg2(40)  <= "111100000111";
  regfileReg2(41)  <= "111100000001";
  regfileReg2(42)  <= "111011111011";
  regfileReg2(43)  <= "111011110101";
  regfileReg2(44)  <= "111011101111";
  regfileReg2(45)  <= "111011101001";
  regfileReg2(46)  <= "111011100011";
  regfileReg2(47)  <= "111011011101";
  regfileReg2(48)  <= "111011010111";
  regfileReg2(49)  <= "111011010001";
  regfileReg2(50)  <= "111011001011";
  regfileReg2(51)  <= "111011000101";
  regfileReg2(52)  <= "111010111111";
  regfileReg2(53)  <= "111010111001";
  regfileReg2(54)  <= "111010110011";
  regfileReg2(55)  <= "111010101101";
  regfileReg2(56)  <= "111010100111";
  regfileReg2(57)  <= "111010100001";
  regfileReg2(58)  <= "111010011011";
  regfileReg2(59)  <= "111010010101";
  regfileReg2(60)  <= "111010001111";
  regfileReg2(61)  <= "111010001010";
  regfileReg2(62)  <= "111010000100";
  regfileReg2(63)  <= "111001111110";
  regfileReg2(64)  <= "111001111000";
  regfileReg2(65)  <= "111001110010";
  regfileReg2(66)  <= "111001101101";
  regfileReg2(67)  <= "111001100111";
  regfileReg2(68)  <= "111001100001";
  regfileReg2(69)  <= "111001011011";
  regfileReg2(70)  <= "111001010110";
  regfileReg2(71)  <= "111001010000";
  regfileReg2(72)  <= "111001001010";
  regfileReg2(73)  <= "111001000101";
  regfileReg2(74)  <= "111000111111";
  regfileReg2(75)  <= "111000111001";
  regfileReg2(76)  <= "111000110100";
  regfileReg2(77)  <= "111000101110";
  regfileReg2(78)  <= "111000101000";
  regfileReg2(79)  <= "111000100011";
  regfileReg2(80)  <= "111000011101";
  regfileReg2(81)  <= "111000011000";
  regfileReg2(82)  <= "111000010010";
  regfileReg2(83)  <= "111000001101";
  regfileReg2(84)  <= "111000000111";
  regfileReg2(85)  <= "111000000010";
  regfileReg2(86)  <= "110111111100";
  regfileReg2(87)  <= "110111110111";
  regfileReg2(88)  <= "110111110010";
  regfileReg2(89)  <= "110111101100";
  regfileReg2(90)  <= "110111100111";
  regfileReg2(91)  <= "110111100001";
  regfileReg2(92)  <= "110111011100";
  regfileReg2(93)  <= "110111010111";
  regfileReg2(94)  <= "110111010010";
  regfileReg2(95)  <= "110111001100";
  regfileReg2(96)  <= "110111000111";
  regfileReg2(97)  <= "110111000010";
  regfileReg2(98)  <= "110110111101";
  regfileReg2(99)  <= "110110111000";
  regfileReg2(100) <= "110110110010";
  regfileReg2(101) <= "110110101101";
  regfileReg2(102) <= "110110101000";
  regfileReg2(103) <= "110110100011";
  regfileReg2(104) <= "110110011110";
  regfileReg2(105) <= "110110011001";
  regfileReg2(106) <= "110110010100";
  regfileReg2(107) <= "110110001111";
  regfileReg2(108) <= "110110001010";
  regfileReg2(109) <= "110110000101";
  regfileReg2(110) <= "110110000000";
  regfileReg2(111) <= "110101111011";
  regfileReg2(112) <= "110101110110";
  regfileReg2(113) <= "110101110010";
  regfileReg2(114) <= "110101101101";
  regfileReg2(115) <= "110101101000";
  regfileReg2(116) <= "110101100011";
  regfileReg2(117) <= "110101011110";
  regfileReg2(118) <= "110101011010";
  regfileReg2(119) <= "110101010101";
  regfileReg2(120) <= "110101010000";
  regfileReg2(121) <= "110101001100";
  regfileReg2(122) <= "110101000111";
  regfileReg2(123) <= "110101000010";
  regfileReg2(124) <= "110100111110";
  regfileReg2(125) <= "110100111001";
  regfileReg2(126) <= "110100110101";
  regfileReg2(127) <= "110100110000";
  regfileReg2(128) <= "110100101100";

end architecture;
